module note_player_tb();

    reg clk, reset, play_enable, generate_next_sample;
    reg [5:0] note_to_load;
    reg [5:0] duration_to_load;
    reg load_new_note;
    wire done_with_note, new_sample_ready, beat;
    wire [15:0] sample_out;

    note_player np(
        .clk(clk),
        .reset(reset),

        .play_enable(play_enable),
        .note_to_load(note_to_load),
        .duration_to_load(duration_to_load),
        .load_new_note(load_new_note),
        .done_with_note(done_with_note),

        .beat(beat),
        .generate_next_sample(generate_next_sample),
        .sample_out(sample_out),
        .new_sample_ready(new_sample_ready)
    );

    beat_generator #(.WIDTH(17), .STOP(1500)) beat_generator(
        .clk(clk),
        .reset(reset),
        .en(1'b1),
        .beat(beat)
    );

    // Clock and reset
    initial begin
        clk = 1'b0;
        reset = 1'b1;
        repeat (4) #5 clk = ~clk;
        reset = 1'b0;
        forever #5 clk = ~clk;
    end

    // Tests
    initial begin
        #33
        play_enable = 1'b1;
        generate_next_sample = 1'b1;
        note_to_load = 6'b000001;
        duration_to_load = 6'd5;
        #10
        $display(sample_out, new_sample_ready, done_with_note);
        
        

    end

//    integer delay;
//    initial begin
//        delay = 2000000;
//        play_enable = 1'b0;
//        load_new_note = 1'b0;
//        @(negedge reset);
//        @(negedge clk);

//        repeat (25) begin
//            @(negedge clk);
//        end 

//        // Start playing
//        $display("Starting playing song 0...");
//        @(negedge clk);
//        play_enable = 1'b1;
//        generate_next_sample = 1'b0;
//        note_to_load = 6'b000001;
//        duration_to_load = 6'd5;
//        load_new_note = 1'b1;
//        @(negedge clk);
//        play_enable = 1'b0;
//        load_new_note = 1'b0;

//        repeat (delay) begin
//            @(negedge clk);
//        end

//        // Pause  
//        $display("Pause...");
//        @(negedge clk);
//        play_enable = 1'b1;
//        @(negedge clk);
//        play_enable = 1'b0;

//        repeat (delay/4) begin
//            @(negedge clk);
//        end
//    end

endmodule
